//-----------------------------------------------------------//
//----------  Configurations Setup for Parameters  ----------//
//-----------------------------------------------------------//
/*
* Description: Change Values of Parameters from this file
*/

package ConfigParams_pkg;
    parameter 	ADDR_WIDTH  =	4;
    parameter   DATA_WIDTH  =   32;
    parameter   CLK_PERIOD  =   10;
endpackage