//-----------------------------------------------------------//
//----------------  Package for all classes  ----------------//
//-----------------------------------------------------------//

package Classes_pkg;
`timescale 1ns/1ps
`include   "TransactionClass.sv"
endpackage